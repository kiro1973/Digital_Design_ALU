`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:05:45 05/18/2021 
// Design Name: 
// Module Name:    OneBitBR 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module OneBitBR(
    input [3:0] OP,
    input A,
    input B,
    input Cin,
    input RES,
    input Cout
    );


endmodule
